	assign sin_table[0] = 40'h0000000000;
	assign sin_table[1] = 40'h0000000996;
	assign sin_table[2] = 40'h000000132A;
	assign sin_table[3] = 40'h0000001CBC;
	assign sin_table[4] = 40'h0000002649;
	assign sin_table[5] = 40'h0000002FD1;
	assign sin_table[6] = 40'h0000003951;
	assign sin_table[7] = 40'h00000042C8;
	assign sin_table[8] = 40'h0000004C35;
	assign sin_table[9] = 40'h0000005596;
	assign sin_table[10] = 40'h0000005EEA;
	assign sin_table[11] = 40'h000000682F;
	assign sin_table[12] = 40'h0000007164;
	assign sin_table[13] = 40'h0000007A88;
	assign sin_table[14] = 40'h0000008398;
	assign sin_table[15] = 40'h0000008C95;
	assign sin_table[16] = 40'h000000957C;
	assign sin_table[17] = 40'h0000009E4C;
	assign sin_table[18] = 40'h000000A703;
	assign sin_table[19] = 40'h000000AFA1;
	assign sin_table[20] = 40'h000000B823;
	assign sin_table[21] = 40'h000000C089;
	assign sin_table[22] = 40'h000000C8D2;
	assign sin_table[23] = 40'h000000D0FB;
	assign sin_table[24] = 40'h000000D905;
	assign sin_table[25] = 40'h000000E0EC;
	assign sin_table[26] = 40'h000000E8B1;
	assign sin_table[27] = 40'h000000F053;
	assign sin_table[28] = 40'h000000F7CF;
	assign sin_table[29] = 40'h000000FF25;
	assign sin_table[30] = 40'h0000010653;
	assign sin_table[31] = 40'h0000010D5A;
	assign sin_table[32] = 40'h0000011436;
	assign sin_table[33] = 40'h0000011AE8;
	assign sin_table[34] = 40'h000001216F;
	assign sin_table[35] = 40'h00000127C8;
	assign sin_table[36] = 40'h0000012DF5;
	assign sin_table[37] = 40'h00000133F2;
	assign sin_table[38] = 40'h00000139C0;
	assign sin_table[39] = 40'h0000013F5E;
	assign sin_table[40] = 40'h00000144CA;
	assign sin_table[41] = 40'h0000014A05;
	assign sin_table[42] = 40'h0000014F0C;
	assign sin_table[43] = 40'h00000153E0;
	assign sin_table[44] = 40'h0000015880;
	assign sin_table[45] = 40'h0000015CEA;
	assign sin_table[46] = 40'h000001611E;
	assign sin_table[47] = 40'h000001651C;
	assign sin_table[48] = 40'h00000168E3;
	assign sin_table[49] = 40'h0000016C73;
	assign sin_table[50] = 40'h0000016FCA;
	assign sin_table[51] = 40'h00000172E8;
	assign sin_table[52] = 40'h00000175CE;
	assign sin_table[53] = 40'h0000017879;
	assign sin_table[54] = 40'h0000017AEB;
	assign sin_table[55] = 40'h0000017D22;
	assign sin_table[56] = 40'h0000017F1E;
	assign sin_table[57] = 40'h00000180DF;
	assign sin_table[58] = 40'h0000018265;
	assign sin_table[59] = 40'h00000183AF;
	assign sin_table[60] = 40'h00000184BE;
	assign sin_table[61] = 40'h0000018591;
	assign sin_table[62] = 40'h0000018627;
	assign sin_table[63] = 40'h0000018681;
	assign sin_table[64] = 40'h00000186A0;
	assign sin_table[65] = 40'h0000018681;
	assign sin_table[66] = 40'h0000018627;
	assign sin_table[67] = 40'h0000018591;
	assign sin_table[68] = 40'h00000184BE;
	assign sin_table[69] = 40'h00000183AF;
	assign sin_table[70] = 40'h0000018265;
	assign sin_table[71] = 40'h00000180DF;
	assign sin_table[72] = 40'h0000017F1E;
	assign sin_table[73] = 40'h0000017D22;
	assign sin_table[74] = 40'h0000017AEB;
	assign sin_table[75] = 40'h0000017879;
	assign sin_table[76] = 40'h00000175CE;
	assign sin_table[77] = 40'h00000172E8;
	assign sin_table[78] = 40'h0000016FCA;
	assign sin_table[79] = 40'h0000016C73;
	assign sin_table[80] = 40'h00000168E3;
	assign sin_table[81] = 40'h000001651C;
	assign sin_table[82] = 40'h000001611E;
	assign sin_table[83] = 40'h0000015CEA;
	assign sin_table[84] = 40'h0000015880;
	assign sin_table[85] = 40'h00000153E0;
	assign sin_table[86] = 40'h0000014F0C;
	assign sin_table[87] = 40'h0000014A05;
	assign sin_table[88] = 40'h00000144CA;
	assign sin_table[89] = 40'h0000013F5E;
	assign sin_table[90] = 40'h00000139C0;
	assign sin_table[91] = 40'h00000133F2;
	assign sin_table[92] = 40'h0000012DF5;
	assign sin_table[93] = 40'h00000127C8;
	assign sin_table[94] = 40'h000001216F;
	assign sin_table[95] = 40'h0000011AE8;
	assign sin_table[96] = 40'h0000011436;
	assign sin_table[97] = 40'h0000010D5A;
	assign sin_table[98] = 40'h0000010653;
	assign sin_table[99] = 40'h000000FF25;
	assign sin_table[100] = 40'h000000F7CF;
	assign sin_table[101] = 40'h000000F053;
	assign sin_table[102] = 40'h000000E8B1;
	assign sin_table[103] = 40'h000000E0EC;
	assign sin_table[104] = 40'h000000D905;
	assign sin_table[105] = 40'h000000D0FB;
	assign sin_table[106] = 40'h000000C8D2;
	assign sin_table[107] = 40'h000000C089;
	assign sin_table[108] = 40'h000000B823;
	assign sin_table[109] = 40'h000000AFA1;
	assign sin_table[110] = 40'h000000A703;
	assign sin_table[111] = 40'h0000009E4C;
	assign sin_table[112] = 40'h000000957C;
	assign sin_table[113] = 40'h0000008C95;
	assign sin_table[114] = 40'h0000008398;
	assign sin_table[115] = 40'h0000007A88;
	assign sin_table[116] = 40'h0000007164;
	assign sin_table[117] = 40'h000000682F;
	assign sin_table[118] = 40'h0000005EEA;
	assign sin_table[119] = 40'h0000005596;
	assign sin_table[120] = 40'h0000004C35;
	assign sin_table[121] = 40'h00000042C8;
	assign sin_table[122] = 40'h0000003951;
	assign sin_table[123] = 40'h0000002FD1;
	assign sin_table[124] = 40'h0000002649;
	assign sin_table[125] = 40'h0000001CBC;
	assign sin_table[126] = 40'h000000132A;
	assign sin_table[127] = 40'h0000000996;
	assign sin_table[128] = 40'h0000000000;
	assign sin_table[129] = 40'hFFFFFFF66A;
	assign sin_table[130] = 40'hFFFFFFECD6;
	assign sin_table[131] = 40'hFFFFFFE344;
	assign sin_table[132] = 40'hFFFFFFD9B7;
	assign sin_table[133] = 40'hFFFFFFD02F;
	assign sin_table[134] = 40'hFFFFFFC6AF;
	assign sin_table[135] = 40'hFFFFFFBD38;
	assign sin_table[136] = 40'hFFFFFFB3CB;
	assign sin_table[137] = 40'hFFFFFFAA6A;
	assign sin_table[138] = 40'hFFFFFFA116;
	assign sin_table[139] = 40'hFFFFFF97D1;
	assign sin_table[140] = 40'hFFFFFF8E9C;
	assign sin_table[141] = 40'hFFFFFF8578;
	assign sin_table[142] = 40'hFFFFFF7C68;
	assign sin_table[143] = 40'hFFFFFF736B;
	assign sin_table[144] = 40'hFFFFFF6A84;
	assign sin_table[145] = 40'hFFFFFF61B4;
	assign sin_table[146] = 40'hFFFFFF58FD;
	assign sin_table[147] = 40'hFFFFFF505F;
	assign sin_table[148] = 40'hFFFFFF47DD;
	assign sin_table[149] = 40'hFFFFFF3F77;
	assign sin_table[150] = 40'hFFFFFF372E;
	assign sin_table[151] = 40'hFFFFFF2F05;
	assign sin_table[152] = 40'hFFFFFF26FB;
	assign sin_table[153] = 40'hFFFFFF1F14;
	assign sin_table[154] = 40'hFFFFFF174F;
	assign sin_table[155] = 40'hFFFFFF0FAD;
	assign sin_table[156] = 40'hFFFFFF0831;
	assign sin_table[157] = 40'hFFFFFF00DB;
	assign sin_table[158] = 40'hFFFFFEF9AD;
	assign sin_table[159] = 40'hFFFFFEF2A6;
	assign sin_table[160] = 40'hFFFFFEEBCA;
	assign sin_table[161] = 40'hFFFFFEE518;
	assign sin_table[162] = 40'hFFFFFEDE91;
	assign sin_table[163] = 40'hFFFFFED838;
	assign sin_table[164] = 40'hFFFFFED20B;
	assign sin_table[165] = 40'hFFFFFECC0E;
	assign sin_table[166] = 40'hFFFFFEC640;
	assign sin_table[167] = 40'hFFFFFEC0A2;
	assign sin_table[168] = 40'hFFFFFEBB36;
	assign sin_table[169] = 40'hFFFFFEB5FB;
	assign sin_table[170] = 40'hFFFFFEB0F4;
	assign sin_table[171] = 40'hFFFFFEAC20;
	assign sin_table[172] = 40'hFFFFFEA780;
	assign sin_table[173] = 40'hFFFFFEA316;
	assign sin_table[174] = 40'hFFFFFE9EE2;
	assign sin_table[175] = 40'hFFFFFE9AE4;
	assign sin_table[176] = 40'hFFFFFE971D;
	assign sin_table[177] = 40'hFFFFFE938D;
	assign sin_table[178] = 40'hFFFFFE9036;
	assign sin_table[179] = 40'hFFFFFE8D18;
	assign sin_table[180] = 40'hFFFFFE8A32;
	assign sin_table[181] = 40'hFFFFFE8787;
	assign sin_table[182] = 40'hFFFFFE8515;
	assign sin_table[183] = 40'hFFFFFE82DE;
	assign sin_table[184] = 40'hFFFFFE80E2;
	assign sin_table[185] = 40'hFFFFFE7F21;
	assign sin_table[186] = 40'hFFFFFE7D9B;
	assign sin_table[187] = 40'hFFFFFE7C51;
	assign sin_table[188] = 40'hFFFFFE7B42;
	assign sin_table[189] = 40'hFFFFFE7A6F;
	assign sin_table[190] = 40'hFFFFFE79D9;
	assign sin_table[191] = 40'hFFFFFE797F;
	assign sin_table[192] = 40'hFFFFFE7960;
	assign sin_table[193] = 40'hFFFFFE797F;
	assign sin_table[194] = 40'hFFFFFE79D9;
	assign sin_table[195] = 40'hFFFFFE7A6F;
	assign sin_table[196] = 40'hFFFFFE7B42;
	assign sin_table[197] = 40'hFFFFFE7C51;
	assign sin_table[198] = 40'hFFFFFE7D9B;
	assign sin_table[199] = 40'hFFFFFE7F21;
	assign sin_table[200] = 40'hFFFFFE80E2;
	assign sin_table[201] = 40'hFFFFFE82DE;
	assign sin_table[202] = 40'hFFFFFE8515;
	assign sin_table[203] = 40'hFFFFFE8787;
	assign sin_table[204] = 40'hFFFFFE8A32;
	assign sin_table[205] = 40'hFFFFFE8D18;
	assign sin_table[206] = 40'hFFFFFE9036;
	assign sin_table[207] = 40'hFFFFFE938D;
	assign sin_table[208] = 40'hFFFFFE971D;
	assign sin_table[209] = 40'hFFFFFE9AE4;
	assign sin_table[210] = 40'hFFFFFE9EE2;
	assign sin_table[211] = 40'hFFFFFEA316;
	assign sin_table[212] = 40'hFFFFFEA780;
	assign sin_table[213] = 40'hFFFFFEAC20;
	assign sin_table[214] = 40'hFFFFFEB0F4;
	assign sin_table[215] = 40'hFFFFFEB5FB;
	assign sin_table[216] = 40'hFFFFFEBB36;
	assign sin_table[217] = 40'hFFFFFEC0A2;
	assign sin_table[218] = 40'hFFFFFEC640;
	assign sin_table[219] = 40'hFFFFFECC0E;
	assign sin_table[220] = 40'hFFFFFED20B;
	assign sin_table[221] = 40'hFFFFFED838;
	assign sin_table[222] = 40'hFFFFFEDE91;
	assign sin_table[223] = 40'hFFFFFEE518;
	assign sin_table[224] = 40'hFFFFFEEBCA;
	assign sin_table[225] = 40'hFFFFFEF2A6;
	assign sin_table[226] = 40'hFFFFFEF9AD;
	assign sin_table[227] = 40'hFFFFFF00DB;
	assign sin_table[228] = 40'hFFFFFF0831;
	assign sin_table[229] = 40'hFFFFFF0FAD;
	assign sin_table[230] = 40'hFFFFFF174F;
	assign sin_table[231] = 40'hFFFFFF1F14;
	assign sin_table[232] = 40'hFFFFFF26FB;
	assign sin_table[233] = 40'hFFFFFF2F05;
	assign sin_table[234] = 40'hFFFFFF372E;
	assign sin_table[235] = 40'hFFFFFF3F77;
	assign sin_table[236] = 40'hFFFFFF47DD;
	assign sin_table[237] = 40'hFFFFFF505F;
	assign sin_table[238] = 40'hFFFFFF58FD;
	assign sin_table[239] = 40'hFFFFFF61B4;
	assign sin_table[240] = 40'hFFFFFF6A84;
	assign sin_table[241] = 40'hFFFFFF736B;
	assign sin_table[242] = 40'hFFFFFF7C68;
	assign sin_table[243] = 40'hFFFFFF8578;
	assign sin_table[244] = 40'hFFFFFF8E9C;
	assign sin_table[245] = 40'hFFFFFF97D1;
	assign sin_table[246] = 40'hFFFFFFA116;
	assign sin_table[247] = 40'hFFFFFFAA6A;
	assign sin_table[248] = 40'hFFFFFFB3CB;
	assign sin_table[249] = 40'hFFFFFFBD38;
	assign sin_table[250] = 40'hFFFFFFC6AF;
	assign sin_table[251] = 40'hFFFFFFD02F;
	assign sin_table[252] = 40'hFFFFFFD9B7;
	assign sin_table[253] = 40'hFFFFFFE344;
	assign sin_table[254] = 40'hFFFFFFECD6;
	assign sin_table[255] = 40'hFFFFFFF66A;
